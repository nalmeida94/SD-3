library verilog;
use verilog.vl_types.all;
entity TB_banco_de_registradores is
end TB_banco_de_registradores;
