library verilog;
use verilog.vl_types.all;
entity TB_extensor_de_sinal is
end TB_extensor_de_sinal;
