library verilog;
use verilog.vl_types.all;
entity TB_pc is
end TB_pc;
