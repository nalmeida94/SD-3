library verilog;
use verilog.vl_types.all;
entity TB_detector_de_flags is
end TB_detector_de_flags;
